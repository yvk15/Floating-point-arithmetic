//This is a PG generator, where P is propagate and G is generate. 
module pg_gen(A, B, P, G);
    input A, B;
    output P, G;

    assign P = A ^ B; 
    assign G = A & B;
endmodule
